//Load a word stored in memory location 120,add 45 to it and stor the
//result in memory location 121

module test_mips32;
  reg clk1, clk2;
  integer k;
  pipe_MIPS32 mips(.clk1(clk1),  .clk2(clk2));
  
  initial begin
    clk1 =0; clk2 =0;
    repeat(20)
      begin
        #5 clk1 = 1; #5 clk2 =0;
        #5 clk1 = 0; #5 clk2 =1;
      end
  end
  
 initial begin
   for(k=0; k<31; k = k+1)
     mips.REG[k] = k;
   mips.MEM[0] = 32'h28010078;  //ADDI R1, R0,120
   mips.MEM[1] = 32'h0ce77800; // OR R7, R7, R7; dummy instn
   mips.MEM[2] = 32'h20220000; //LW R2, 0(R1)
   mips.MEM[3] = 32'h0ce77800; // OR R7, R7, R7; dummy instn
   mips.MEM[4] = 32'h2842002d; //ADDI R2,R2 45
   mips.MEM[5] = 32'h0ce77800; // OR R7, R7, R7; dummy instn
   mips.MEM[6] = 32'h24220001; //SW R2, 1(R1)
   mips.MEM[7] = 32'hfc000000; //hlt
   
   mips.MEM[120] = 85;
   
  mips.HALTED = 0;
  mips.PC = 0;
  mips. TAKEN_BRANCH =0;
   
   #500 $display ("MEM[120]: %4d\n MEM[121] : %4d", mips.MEM[120], mips.MEM[121]);
 end
  
  
   initial 
     begin
       $dumpfile("waveform.vcd");
     $dumpvars(0,test_mips32);
     end
   

    initial begin
     #600 $finish;
   end
 
   endmodule
   